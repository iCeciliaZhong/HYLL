`define MATRIX_SIZE   16
`define COLOR_DEPTH   8
`define ADDR_WIDTH    8

