`define MATRIX_SIZE   8
`define COLOR_DEPTH   8
`define ADDR_WIDTH    6
//`define ILA 